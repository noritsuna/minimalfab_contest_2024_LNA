* Created by KLayout

* cell base_Rev0.94
.SUBCKT base_Rev0.94
* device instance $1 r0 *1 204,-439.5 NMOS
M$1 5 9 1 1 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $2 r0 *1 204,-599.5 NMOS
M$2 5 7 8 8 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $3 r0 *1 44,-439.5 NMOS
M$3 91 89 90 90 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $4 r0 *1 44,-599.5 NMOS
M$4 8 3 6 6 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $5 r0 *1 -436,-439.5 NMOS
M$5 70 67 25 25 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $6 r0 *1 -436,-599.5 NMOS
M$6 6 3 3 3 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $7 r0 *1 -596,-439.5 NMOS
M$7 94 92 93 93 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $8 r0 *1 -596,-599.5 NMOS
M$8 73 76 86 86 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $9 r0 *1 204,200.5 NMOS
M$9 68 65 23 23 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $10 r0 *1 204,40.5 NMOS
M$10 87 82 77 77 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $11 r0 *1 44,200.5 NMOS
M$11 97 95 96 96 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $12 r0 *1 44,40.5 NMOS
M$12 71 74 84 84 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $13 r0 *1 -436,200.5 NMOS
M$13 69 66 24 24 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $14 r0 *1 -436,40.5 NMOS
M$14 88 83 78 78 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $15 r0 *1 -596,200.5 NMOS
M$15 100 98 99 99 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $16 r0 *1 -596,40.5 NMOS
M$16 72 75 85 85 NMOS L=10U W=10U AS=229P AD=229P PS=64U PD=64U
* device instance $24 r0 *1 356.5,-442 PRES
R$24 9 4 28800 PRES
* device instance $25 r0 *1 -43.5,-362 PRES
R$25 52 46 3600 PRES
* device instance $26 r0 *1 -43.5,-442 PRES
R$26 81 55 3600 PRES
* device instance $27 r0 *1 -123.5,-362 PRES
R$27 40 49 3600 PRES
* device instance $28 r0 *1 -123.5,-442 PRES
R$28 58 43 3600 PRES
* device instance $29 r0 *1 -203.5,-362 PRES
R$29 34 28 3600 PRES
* device instance $30 r0 *1 -203.5,-442 PRES
R$30 61 37 3600 PRES
* device instance $31 r0 *1 -283.5,-362 PRES
R$31 19 31 3600 PRES
* device instance $32 r0 *1 -283.5,-442 PRES
R$32 64 22 3600 PRES
* device instance $33 r0 *1 596.5,278 PRES
R$33 50 44 3600 PRES
* device instance $34 r0 *1 596.5,198 PRES
R$34 79 53 3600 PRES
* device instance $35 r0 *1 516.5,278 PRES
R$35 38 47 3600 PRES
* device instance $36 r0 *1 516.5,198 PRES
R$36 56 41 3600 PRES
* device instance $37 r0 *1 436.5,278 PRES
R$37 32 26 3600 PRES
* device instance $38 r0 *1 436.5,198 PRES
R$38 59 35 3600 PRES
* device instance $39 r0 *1 356.5,278 PRES
R$39 17 29 3600 PRES
* device instance $40 r0 *1 356.5,198 PRES
R$40 62 20 3600 PRES
* device instance $41 r0 *1 -43.5,278 PRES
R$41 51 45 3600 PRES
* device instance $42 r0 *1 -43.5,198 PRES
R$42 80 54 3600 PRES
* device instance $43 r0 *1 -123.5,278 PRES
R$43 39 48 3600 PRES
* device instance $44 r0 *1 -123.5,198 PRES
R$44 57 42 3600 PRES
* device instance $45 r0 *1 -203.5,278 PRES
R$45 33 27 3600 PRES
* device instance $46 r0 *1 -203.5,198 PRES
R$46 60 36 3600 PRES
* device instance $47 r0 *1 -283.5,278 PRES
R$47 18 30 3600 PRES
* device instance $48 r0 *1 -283.5,198 PRES
R$48 63 21 3600 PRES
* device instance $49 r0 *1 559.75,-98.5 TINCAP
C$49 8 9 1.656e-12 TINCAP
.ENDS base_Rev0.94
